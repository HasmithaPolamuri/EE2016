module carry(c, a,b);

input a;
input b;
output c;

and(c,a,b);



endmodule
